//对汇编码的修改包括：32位立即数相关，几处笔误，blt改为bltz，Exception后添加返回（此处及中断是否应该返回的是26号而非31号？）
module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	localparam ROM_SIZE = 128;
	(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

	integer i;
	initial begin
		ROMDATA[0]<=32'b00001000000000000000000000000011;	//j Main
		ROMDATA[1]<=32'b00001000000000000000000001001011;	//j Interruption
		ROMDATA[2]<=32'b00001000000000000000000001010000;	//j Exception
		ROMDATA[3]<=32'b00100000000111010000000000000000;	//Main:    addi $sp,$zero,0
		ROMDATA[4]<=32'b00111100000010000100000000000000;	//lui $t0,16384
		ROMDATA[5]<=32'b10101101000000000000000000001000;	//sw $zero,8($t0)
		ROMDATA[6]<=32'b00111100000010011000100010001000;	//lui $t1,34952
		ROMDATA[7]<=32'b00100001001010011000100010001000;	//addi $t1,$t1,34952
		ROMDATA[8]<=32'b10101101000010010000000000000000;	//sw $t1,0($t0)
		ROMDATA[9]<=32'b00111100000010011111111111111111;	//lui $t1,65535
		ROMDATA[10]<=32'b00100001001010011111111111111111;	//addi $t1,$t1,65535
		ROMDATA[11]<=32'b10101101000010010000000000000100;	//sw $t1,4($t0)		
		ROMDATA[12]<=32'b00100000000010010000000000000011;	//addi $t1,$zero,3
		ROMDATA[13]<=32'b10101101000010010000000000001000;	//sw $t1,8($t0)
		ROMDATA[14]<=32'b00100000000010010000000000000011;	//addi $t1,$zero,3
		ROMDATA[15]<=32'b10101101000010010000000000100000;	//sw $t1,32($t0)
		ROMDATA[16]<=32'b10001101000010010000000000100000;	//load_number1:    lw $t1,32($t0) 	
		ROMDATA[17]<=32'b00110001001010100000000000001000;	//andi $t2,$t1,8		 
		ROMDATA[18]<=32'b00010000000010101111111111111101;	//beq $t2,$zero,load_number1 
		ROMDATA[19]<=32'b10001101000100000000000000011100;	//lw $s0,28($t0)		
		ROMDATA[20]<=32'b10001101000010010000000000100000;	//load_number2:    lw $t1,32($t0)
		ROMDATA[21]<=32'b00110001001010100000000000001000;	//andi $t2,$t1,8
		ROMDATA[22]<=32'b00010000000010101111111111111101;	//beq $t2,$zero,load_number2
		ROMDATA[23]<=32'b10001101000100010000000000011100;	//lw $s1,28($t0)		
		ROMDATA[24]<=32'b00111100000011000011111111111111;	//lui $t4,16383
		ROMDATA[25]<=32'b00100001100011001111110000000000;	//addi $t4,$t4,64512
		ROMDATA[26]<=32'b00000010000011000100100000100000;	//add $t1,$s0,$t4
		ROMDATA[27]<=32'b10001101001100100000000000000000;	//lw $s2,0($t1)
		ROMDATA[28]<=32'b00000010001011000100100000100000;	//add $t1,$s1,$t4
		ROMDATA[29]<=32'b10001101001100110000000000000000;	//lw $s3,0($t1)
		ROMDATA[30]<=32'b00000010000000000010000000100000;	//add $a0,$s0,$zero
		ROMDATA[31]<=32'b00000010001000000010100000100000;	//add $a1,$s1,$zero
		ROMDATA[32]<=32'b00010000101001000000000000000111;	//compare:    beq $a0,$a1,exit
		ROMDATA[33]<=32'b00000000101001000110000000100010;	//sub $t4,$a1,$a0
		ROMDATA[34]<=32'b01001001100000000000000000000011;	//bltz $t4,minus
		ROMDATA[35]<=32'b00000000100000000100100000100000;	//add $t1,$a0,$zero
		ROMDATA[36]<=32'b00000000101000000010000000100000;	//add $a0,$a1,$zero
		ROMDATA[37]<=32'b00000001000000000010100000100000;	//add $a1,$t0,$zero
		ROMDATA[38]<=32'b00000000100001010010000000100010;	//minus:    sub $a0,$a0,$a1
		ROMDATA[39]<=32'b00001000000000000000000000100000;	//j compare
		ROMDATA[40]<=32'b10001101000010010000000000100000;	//exit:    lw $t1,32($t0) 	
		ROMDATA[41]<=32'b00110001001010100000000000000100;	//andi $t2,$t1,4		 
		ROMDATA[42]<=32'b00010000000010101111111111111101;	//beq $t2,$zero,exit
		ROMDATA[43]<=32'b10101101000001000000000000011000;	//sw $a0,24($t0)
		ROMDATA[44]<=32'b10101101000001000000000000001100;	//display_result:    sw $a0,12($t0)
		ROMDATA[45]<=32'b00000000000100100101011001000000;	//decode1:    sll $t2,$s2,25
		ROMDATA[46]<=32'b00000000000010100101011001000010;	//srl $t2,$t2,25
		ROMDATA[47]<=32'b00000000000100110101111001000000;	//sll $t3,$s3,25
		ROMDATA[48]<=32'b00000000000010110101101110000010;	//srl $t3,$t3,14
		ROMDATA[49]<=32'b00100001010010100000000010000000;	//addi $t2,$t2,128
		ROMDATA[50]<=32'b00000001010010110101000000100000;	//add $t2,$t2,$t3
		ROMDATA[51]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)
		ROMDATA[52]<=32'b00001100000000000000000001001011;	//jal Interruption
		ROMDATA[53]<=32'b00000000000100100101010010000000;	//decode2:    sll $t2,$s2,18
		ROMDATA[54]<=32'b00000000000010100101011001000010;	//srl $t2,$t2,25
		ROMDATA[55]<=32'b00000000000100110101110010000000;	//sll $t3,$s3,18
		ROMDATA[56]<=32'b00000000000010110101111001000010;	//srl $t3,$t3,25
		ROMDATA[57]<=32'b00000000000010110101101011000000;	//sll $t3,$t3,11
		ROMDATA[58]<=32'b00100001010010100000000100000000;	//addi $t2,$t2,256
		ROMDATA[59]<=32'b00000001010010110101000000100000;	//add $t2,$t2,$t3
		ROMDATA[60]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)
		ROMDATA[61]<=32'b00001100000000000000000001001011;	//jal Interruption
		ROMDATA[62]<=32'b00000000000100100101001011000000;	//decode3:    sll $t2,$s2,11
		ROMDATA[63]<=32'b00000000000010100101011001000010;	//srl $t2,$t2,25
		ROMDATA[64]<=32'b00000000000100110101101011000000;	//sll $t3,$s3,11
		ROMDATA[65]<=32'b00000000000010110101111001000010;	//srl $t3,$t3,25
		ROMDATA[66]<=32'b00000000000010110101101011000000;	//sll $t3,$t3,11
		ROMDATA[67]<=32'b00100001010010100000001000000000;	//addi $t2,$t2,512
		ROMDATA[68]<=32'b00000001010010110101000000100000;	//add $t2,$t2,$t3
		ROMDATA[69]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)
		ROMDATA[70]<=32'b00001100000000000000000001001011;	//jal Interruption
		ROMDATA[71]<=32'b00100000000010100000010000000000;	//decode4:    addi $t2,$zero,1024
		ROMDATA[72]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)
		ROMDATA[73]<=32'b00001100000000000000000001001011;	//jal Interruption
		ROMDATA[74]<=32'b00001100000000000000000000101101;	//jal decode1
		ROMDATA[75]<=32'b10001101000010010000000000001000;	//Interruption:    lw $t1,8($t0)
		ROMDATA[76]<=32'b00100000000010010000000000000001;	//addi $t1,$zero,1
		ROMDATA[77]<=32'b10101101000010010000000000001000;	//sw $t1,8($t0)
		ROMDATA[78]<=32'b00000000000000000000000000000000;	//sll $zero,$zero,0
		ROMDATA[79]<=32'b00000011111000000000000000001000;	//jr $ra
		ROMDATA[80]<=32'b00000000000000000000000000000000;	//Exception:    sll $zero,$zero,0
	    for (i=81;i<ROM_SIZE;i=i+1) begin
            ROMDATA[i] <= 32'b0;
        end
	end
	
	always@(*) Instruction<=(Address[9:2] < ROM_SIZE)?ROMDATA[Address[9:2]]:32'b0;
	
endmodule
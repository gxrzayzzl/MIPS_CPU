//对汇编码的修改包括：32位立即数相关，几处笔误，blt改为bltz，Exception后添加返回（此处及中断是否应该返回的是26号而非31号？）
module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	localparam ROM_SIZE = 128;
	(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

	integer i;
	initial begin
		ROMDATA[0]<=32'b00001000000000000000000000000011;	//j Main
		ROMDATA[1]<=32'b00001000000000000000000001001100;	//j Interruption
		ROMDATA[2]<=32'b00001000000000000000000001010011;	//j Exception
		ROMDATA[3]<=32'b00100000000111010000000000000000;	//Main:    addi $sp,$zero,0 c
		ROMDATA[4]<=32'b00111100000010000100000000000000;	//lui $t0,16384             10
		ROMDATA[5]<=32'b10101101000000000000000000001000;	//sw $zero,8($t0)           14
		ROMDATA[6]<=32'b00111100000010011111111111111111;	//lui $t1,65535             18
		ROMDATA[7]<=32'b10101101000010010000000000000000;	//ori $t1,$t1,60000         1c
		ROMDATA[8]<=32'b10101101000010010000000000000000;	//sw $t1,0($t0)             20
		ROMDATA[9]<=32'b00111100000010011111111111111111;	//lui $t1,65535             24
		ROMDATA[10]<=32'b00100001001010011111111111111111;	//addi $t1,$t1,65535        28
		ROMDATA[11]<=32'b10101101000010010000000000000100;	//sw $t1,4($t0)		        2c
		ROMDATA[12]<=32'b00100000000010010000000000000010;	//addi $t1,$zero,2          30
		ROMDATA[13]<=32'b10101101000010010000000000001000;	//sw $t1,8($t0)             34
		ROMDATA[14]<=32'b00100000000010010000000000000011;	//addi $t1,$zero,3          38
		ROMDATA[15]<=32'b10101101000010010000000000100000;	//sw $t1,32($t0)            3c
		ROMDATA[16]<=32'b10001101000010010000000000100000;	//load_number1:    lw $t1,32($t0) 40	
		ROMDATA[17]<=32'b00110001001010100000000000001000;	//andi $t2,$t1,8		 
		ROMDATA[18]<=32'b00010000000010101111111111111101;	//beq $t2,$zero,load_number1 
		ROMDATA[19]<=32'b10001101000100000000000000011100;	//lw $s0,28($t0)		
		ROMDATA[20]<=32'b10001101000010010000000000100000;	//load_number2:    lw $t1,32($t0) 50
		ROMDATA[21]<=32'b00110001001010100000000000001000;	//andi $t2,$t1,8                  54
		ROMDATA[22]<=32'b00010000000010101111111111111101;	//beq $t2,$zero,load_number2      58
		ROMDATA[23]<=32'b10001101000100010000000000011100;	//lw $s1,28($t0)                  5c
		ROMDATA[24]<=32'b00100000000011000000010000000000;	//addi $t4,$zero,1024             60
		ROMDATA[25]<=32'b00000000000100000100100010000000;	//sll $t1,$s0,2                   64
		ROMDATA[26]<=32'b00000001001011000100100000100000;	//add $t1,$t1,$t4                 68
		ROMDATA[27]<=32'b10001101001100100000000000000000;	//lw $s2,0($t1)                   6c
		ROMDATA[28]<=32'b00000000000100010100100010000000;	//sll $t1,$s1,2                   70
		ROMDATA[29]<=32'b00000001001011000100100000100000;	//add $t1,$t1,$t4                 74
		ROMDATA[30]<=32'b10001101001100110000000000000000;	//lw $s3,0($t1)                   78
		ROMDATA[31]<=32'b00000010000000000010000000100000;	//add $a0,$s0,$zero
		ROMDATA[32]<=32'b00000010001000000010100000100000;	//add $a1,$s1,$zero
		ROMDATA[33]<=32'b00010000101001000000000000000111;	//compare:    beq $a0,$a1,exit
		ROMDATA[34]<=32'b00000000101001000110000000100010;	//sub $t4,$a1,$a0
		ROMDATA[35]<=32'b00000101100000000000000000000011;	//bltz $t4,minus
		ROMDATA[36]<=32'b00000000100000000100100000100000;	//add $t1,$a0,$zero
		ROMDATA[37]<=32'b00000000101000000010000000100000;	//add $a0,$a1,$zero
		ROMDATA[38]<=32'b00000001001000000010100000100000;	//add $a1,$t1,$zero         
		ROMDATA[39]<=32'b00000000100001010010000000100010;	//minus:    sub $a0,$a0,$a1 9c
		ROMDATA[40]<=32'b00001000000000000000000000100001;	//j compare                 a0
		ROMDATA[41]<=32'b10001101000010010000000000100000;	//exit:    lw $t1,32($t0)   a4	
		ROMDATA[42]<=32'b00110001001010100000000000000110;	//andi $t2,$t1,4		    a8
		ROMDATA[43]<=32'b00010000000010101111111111111101;	//beq $t2,$zero,exit        ac
		ROMDATA[44]<=32'b10101101000001000000000000011000;	//sw $a0,24($t0)            b0
		ROMDATA[45]<=32'b10101101000001000000000000001100;	//display_result:    sw $a0,12($t0)  b4
		ROMDATA[46]<=32'b00000000000100100101011001000000;	//decode1:    sll $t2,$s2,25         b8
		ROMDATA[47]<=32'b00000000000010100101011001000010;	//srl $t2,$t2,25                     bc
		ROMDATA[48]<=32'b00000000000100110101111001000000;	//sll $t3,$s3,25                     c0
		ROMDATA[49]<=32'b00000000000010110101101110000010;	//srl $t3,$t3,14                     c4
		ROMDATA[50]<=32'b00100001010010100000000010000000;	//addi $t2,$t2,128                   c8
		ROMDATA[51]<=32'b00000001010010110101000000100000;	//add $t2,$t2,$t3                    cc
		ROMDATA[52]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)                     d0
		ROMDATA[53]<=32'b00001100000000000000000001001100;	//jal Interruption                   d4
		ROMDATA[54]<=32'b00000000000100100101010010000000;	//decode2:    sll $t2,$s2,18         d8
		ROMDATA[55]<=32'b00000000000010100101011001000010;	//srl $t2,$t2,25                     dc
		ROMDATA[56]<=32'b00000000000100110101110010000000;	//sll $t3,$s3,18                     e0
		ROMDATA[57]<=32'b00000000000010110101111001000010;	//srl $t3,$t3,25                     e4  
		ROMDATA[58]<=32'b00000000000010110101101011000000;	//sll $t3,$t3,11                     e8
		ROMDATA[59]<=32'b00100001010010100000000100000000;	//addi $t2,$t2,256                   ec
		ROMDATA[60]<=32'b00000001010010110101000000100000;	//add $t2,$t2,$t3                    f0 
		ROMDATA[61]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)                     f4
		ROMDATA[62]<=32'b00001100000000000000000001001100;	//jal Interruption                   f8
		ROMDATA[63]<=32'b00000000000100100101001011000000;	//decode3:    sll $t2,$s2,11         fc
		ROMDATA[64]<=32'b00000000000010100101011001000010;	//srl $t2,$t2,25                     100
		ROMDATA[65]<=32'b00000000000100110101101011000000;	//sll $t3,$s3,11                     104
		ROMDATA[66]<=32'b00000000000010110101111001000010;	//srl $t3,$t3,25                     108
		ROMDATA[67]<=32'b00000000000010110101101011000000;	//sll $t3,$t3,11                     10c
		ROMDATA[68]<=32'b00100001010010100000001000000000;	//addi $t2,$t2,512                   110
		ROMDATA[69]<=32'b00000001010010110101000000100000;	//add $t2,$t2,$t3                    114
		ROMDATA[70]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)                     118
		ROMDATA[71]<=32'b00001100000000000000000001001100;	//jal Interruption                   11c
		ROMDATA[72]<=32'b00100000000010100000010000000000;	//decode4:    addi $t2,$zero,1024    120
 		ROMDATA[73]<=32'b10101101000010100000000000010100;	//sw $t2,20($t0)                     124
		ROMDATA[74]<=32'b00001100000000000000000001001100;	//jal Interruption                   128
		ROMDATA[75]<=32'b00001100000000000000000000101110;	//jal decode1                        12c
		ROMDATA[76]<=32'b10001101000010010000000000001000;	//Interruption:    lw $t1,8($t0)     130
		ROMDATA[77]<=32'b00100000000010010000000000000011;	//addi $t1,$zero,3                   134
		ROMDATA[78]<=32'b10101101000010010000000000001000;	//sw $t1,8($t0)                      138
		ROMDATA[79]<=32'b00000000000000000000000000000000;	//sll $zero,$zero,0                  13c
		ROMDATA[80]<=32'b00100000000010010000000000000010;	//addi $t1,$zero,2                   140
		ROMDATA[81]<=32'b10101101000010010000000000001000;	//sw $t1,8($t0)                      144
		ROMDATA[82]<=32'b00000011111000000000000000001000;	//jr $ra                             148
		ROMDATA[83]<=32'b00000000000000000000000000000000;	//Exception:    nop
		ROMDATA[84]<=32'b00001000000000000000000001010011;	//j Exception
	    for (i=85;i<ROM_SIZE;i=i+1) begin
            ROMDATA[i] <= 32'b0;
        end
	end
	
	always@(*) Instruction<=(Address[9:2] < ROM_SIZE)?ROMDATA[Address[9:2]]:32'b0;
	
endmodule
module DataMemory(
input reset,
input sysclk,
input clk,
input Uart_Rx,
input read_enable,
input write_enable,
input[31:0] address,
input[31:0] writedata,
input[7:0] switch,
output[7:0] led,
output[17:0] tube,
output Uart_Tx,
output wire[31:0] readdata,
output if_continue
    );
    
reg[31:0] memory[255:0];
reg[31:0] tmp;
assign readdata = tmp;
reg[17:0] tubereg;
assign tube = tubereg;
reg[7:0] ledreg;
assign led = ledreg;
reg[7:0] UartWriteData;
wire[7:0] UartReadData;

reg[31:0] timer_TH;
wire[31:0] timer_TL;
reg[1:0] timer_CON_W;
wire timer_CON_R;
reg[1:0] Uart_CON_W;
wire[2:0] Uart_CON_R;

reg Uart_send_trigger;
reg Uart_state_trigger;

integer i;

    always@ (*)
    if(read_enable && address == 32'h40000020) Uart_state_trigger = 1'b1;
    else Uart_state_trigger = 1'b0;

    always@ (*)
    if(read_enable) begin
            case(address)   
                32'h4000001c : tmp = {24'b0,UartReadData};
                32'h40000010 : tmp = {24'b0,switch};
                32'h40000020 : tmp = {27'b0,Uart_CON_R,Uart_CON_W};
                32'h40000008 : tmp = {29'b0,timer_CON_R,timer_CON_W};
                32'h40000004 : tmp = timer_TL;
                32'd1024 :tmp = {11'b0,21'b011111101111110111111};
                32'd1028 :tmp = {11'b0,21'b011111101111110000110};
                32'd1032 :tmp = {11'b0,21'b011111101111111011011};
                32'd1036 :tmp = {11'b0,21'b011111101111111001111};
                32'd1040 :tmp = {11'b0,21'b011111101111111100110};
                32'd1044 :tmp = {11'b0,21'b011111101111111101101};
                32'd1048 :tmp = {11'b0,21'b011111101111111111101};
                32'd1052 :tmp = {11'b0,21'b011111101111110000111};
                32'd1056 :tmp = {11'b0,21'b011111101111111111111};
                32'd1060 :tmp = {11'b0,21'b011111101111111101111};
                32'd1064 :tmp = {11'b0,21'b011111100001100111111};
                32'd1068 :tmp = {11'b0,21'b011111100001100000110};
                32'd1072 :tmp = {11'b0,21'b011111100001101011011};
                32'd1076 :tmp = {11'b0,21'b011111100001101001111};
                32'd1080 :tmp = {11'b0,21'b011111100001101100110};
                32'd1084 :tmp = {11'b0,21'b011111100001101101101};
                32'd1088 :tmp = {11'b0,21'b011111100001101111101};
                32'd1092 :tmp = {11'b0,21'b011111100001100000111};
                32'd1096 :tmp = {11'b0,21'b011111100001101111111};
                32'd1100 :tmp = {11'b0,21'b011111100001101101111};
                32'd1104 :tmp = {11'b0,21'b011111110110110111111};
                32'd1108 :tmp = {11'b0,21'b011111110110110000110};
                32'd1112 :tmp = {11'b0,21'b011111110110111011011};
                32'd1116 :tmp = {11'b0,21'b011111110110111001111};
                32'd1120 :tmp = {11'b0,21'b011111110110111100110};
                32'd1124 :tmp = {11'b0,21'b011111110110111101101};
                32'd1128 :tmp = {11'b0,21'b011111110110111111101};
                32'd1132 :tmp = {11'b0,21'b011111110110110000111};
                32'd1136 :tmp = {11'b0,21'b011111110110111111111};
                32'd1140 :tmp = {11'b0,21'b011111110110111101111};
                32'd1144 :tmp = {11'b0,21'b011111110011110111111};
                32'd1148 :tmp = {11'b0,21'b011111110011110000110};
                32'd1152 :tmp = {11'b0,21'b011111110011111011011};
                32'd1156 :tmp = {11'b0,21'b011111110011111001111};
                32'd1160 :tmp = {11'b0,21'b011111110011111100110};
                32'd1164 :tmp = {11'b0,21'b011111110011111101101};
                32'd1168 :tmp = {11'b0,21'b011111110011111111101};
                32'd1172 :tmp = {11'b0,21'b011111110011110000111};
                32'd1176 :tmp = {11'b0,21'b011111110011111111111};
                32'd1180 :tmp = {11'b0,21'b011111110011111101111};
                32'd1184 :tmp = {11'b0,21'b011111111001100111111};
                32'd1188 :tmp = {11'b0,21'b011111111001100000110};
                32'd1192 :tmp = {11'b0,21'b011111111001101011011};
                32'd1196 :tmp = {11'b0,21'b011111111001101001111};
                32'd1200 :tmp = {11'b0,21'b011111111001101100110};
                32'd1204 :tmp = {11'b0,21'b011111111001101101101};
                32'd1208 :tmp = {11'b0,21'b011111111001101111101};
                32'd1212 :tmp = {11'b0,21'b011111111001100000111};
                32'd1216 :tmp = {11'b0,21'b011111111001101111111};
                32'd1220 :tmp = {11'b0,21'b011111111001101101111};
                32'd1224 :tmp = {11'b0,21'b011111111011010111111};
                32'd1228 :tmp = {11'b0,21'b011111111011010000110};
                32'd1232 :tmp = {11'b0,21'b011111111011011011011};
                32'd1236 :tmp = {11'b0,21'b011111111011011001111};
                32'd1240 :tmp = {11'b0,21'b011111111011011100110};
                32'd1244 :tmp = {11'b0,21'b011111111011011101101};
                32'd1248 :tmp = {11'b0,21'b011111111011011111101};
                32'd1252 :tmp = {11'b0,21'b011111111011010000111};
                32'd1256 :tmp = {11'b0,21'b011111111011011111111};
                32'd1260 :tmp = {11'b0,21'b011111111011011101111};
                32'd1264 :tmp = {11'b0,21'b011111111111010111111};
                32'd1268 :tmp = {11'b0,21'b011111111111010000110};
                32'd1272 :tmp = {11'b0,21'b011111111111011011011};
                32'd1276 :tmp = {11'b0,21'b011111111111011001111};
                32'd1280 :tmp = {11'b0,21'b011111111111011100110};
                32'd1284 :tmp = {11'b0,21'b011111111111011101101};
                32'd1288 :tmp = {11'b0,21'b011111111111011111101};
                32'd1292 :tmp = {11'b0,21'b011111111111010000111};
                32'd1296 :tmp = {11'b0,21'b011111111111011111111};
                32'd1300 :tmp = {11'b0,21'b011111111111011101111};
                32'd1304 :tmp = {11'b0,21'b011111100001110111111};
                32'd1308 :tmp = {11'b0,21'b011111100001110000110};
                32'd1312 :tmp = {11'b0,21'b011111100001111011011};
                32'd1316 :tmp = {11'b0,21'b011111100001111001111};
                32'd1320 :tmp = {11'b0,21'b011111100001111100110};
                32'd1324 :tmp = {11'b0,21'b011111100001111101101};
                32'd1328 :tmp = {11'b0,21'b011111100001111111101};
                32'd1332 :tmp = {11'b0,21'b011111100001110000111};
                32'd1336 :tmp = {11'b0,21'b011111100001111111111};
                32'd1340 :tmp = {11'b0,21'b011111100001111101111};
                32'd1344 :tmp = {11'b0,21'b011111111111110111111};
                32'd1348 :tmp = {11'b0,21'b011111111111110000110};
                32'd1352 :tmp = {11'b0,21'b011111111111111011011};
                32'd1356 :tmp = {11'b0,21'b011111111111111001111};
                32'd1360 :tmp = {11'b0,21'b011111111111111100110};
                32'd1364 :tmp = {11'b0,21'b011111111111111101101};
                32'd1368 :tmp = {11'b0,21'b011111111111111111101};
                32'd1372 :tmp = {11'b0,21'b011111111111110000111};
                32'd1376 :tmp = {11'b0,21'b011111111111111111111};
                32'd1380 :tmp = {11'b0,21'b011111111111111101111};
                32'd1384 :tmp = {11'b0,21'b011111111011110111111};
                32'd1388 :tmp = {11'b0,21'b011111111011110000110};
                32'd1392 :tmp = {11'b0,21'b011111111011111011011};
                32'd1396 :tmp = {11'b0,21'b011111111011111001111};
                32'd1400 :tmp = {11'b0,21'b011111111011111100110};
                32'd1404 :tmp = {11'b0,21'b011111111011111101101};
                32'd1408 :tmp = {11'b0,21'b011111111011111111101};
                32'd1412 :tmp = {11'b0,21'b011111111011110000111};
                32'd1416 :tmp = {11'b0,21'b011111111011111111111};
                32'd1420 :tmp = {11'b0,21'b011111111011111101111};
                32'd1424 :tmp = {11'b0,21'b000011001111110111111};
                32'd1428 :tmp = {11'b0,21'b000011001111110000110};
                32'd1432 :tmp = {11'b0,21'b000011001111111011011};
                32'd1436 :tmp = {11'b0,21'b000011001111111001111};
                32'd1440 :tmp = {11'b0,21'b000011001111111100110};
                32'd1444 :tmp = {11'b0,21'b000011001111111101101};
                32'd1448 :tmp = {11'b0,21'b000011001111111111101};
                32'd1452 :tmp = {11'b0,21'b000011001111110000111};
                32'd1456 :tmp = {11'b0,21'b000011001111111111111};
                32'd1460 :tmp = {11'b0,21'b000011001111111101111};
                32'd1464 :tmp = {11'b0,21'b000011000001100111111};
                32'd1468 :tmp = {11'b0,21'b000011000001100000110};
                32'd1472 :tmp = {11'b0,21'b000011000001101011011};
                32'd1476 :tmp = {11'b0,21'b000011000001101001111};
                32'd1480 :tmp = {11'b0,21'b000011000001101100110};
                32'd1484 :tmp = {11'b0,21'b000011000001101101101};
                32'd1488 :tmp = {11'b0,21'b000011000001101111101};
                32'd1492 :tmp = {11'b0,21'b000011000001100000111};
                32'd1496 :tmp = {11'b0,21'b000011000001101111111};
                32'd1500 :tmp = {11'b0,21'b000011000001101101111};
                32'd1504 :tmp = {11'b0,21'b000011010110110111111};
                32'd1508 :tmp = {11'b0,21'b000011010110110000110};
                32'd1512 :tmp = {11'b0,21'b000011010110111011011};
                32'd1516 :tmp = {11'b0,21'b000011010110111001111};
                32'd1520 :tmp = {11'b0,21'b000011010110111100110};
                32'd1524 :tmp = {11'b0,21'b000011010110111101101};
                32'd1528 :tmp = {11'b0,21'b000011010110111111101};
                32'd1532 :tmp = {11'b0,21'b000011010110110000111};
                32'd1536 :tmp = {11'b0,21'b000011010110111111111};
                32'd1540 :tmp = {11'b0,21'b000011010110111101111};
                32'd1544 :tmp = {11'b0,21'b000011010011110111111};
                32'd1548 :tmp = {11'b0,21'b000011010011110000110};
                32'd1552 :tmp = {11'b0,21'b000011010011111011011};
                32'd1556 :tmp = {11'b0,21'b000011010011111001111};
                32'd1560 :tmp = {11'b0,21'b000011010011111100110};
                32'd1564 :tmp = {11'b0,21'b000011010011111101101};
                32'd1568 :tmp = {11'b0,21'b000011010011111111101};
                32'd1572 :tmp = {11'b0,21'b000011010011110000111};
                32'd1576 :tmp = {11'b0,21'b000011010011111111111};
                32'd1580 :tmp = {11'b0,21'b000011010011111101111};
                32'd1584 :tmp = {11'b0,21'b000011011001100111111};
                32'd1588 :tmp = {11'b0,21'b000011011001100000110};
                32'd1592 :tmp = {11'b0,21'b000011011001101011011};
                32'd1596 :tmp = {11'b0,21'b000011011001101001111};
                32'd1600 :tmp = {11'b0,21'b000011011001101100110};
                32'd1604 :tmp = {11'b0,21'b000011011001101101101};
                32'd1608 :tmp = {11'b0,21'b000011011001101111101};
                32'd1612 :tmp = {11'b0,21'b000011011001100000111};
                32'd1616 :tmp = {11'b0,21'b000011011001101111111};
                32'd1620 :tmp = {11'b0,21'b000011011001101101111};
                32'd1624 :tmp = {11'b0,21'b000011011011010111111};
                32'd1628 :tmp = {11'b0,21'b000011011011010000110};
                32'd1632 :tmp = {11'b0,21'b000011011011011011011};
                32'd1636 :tmp = {11'b0,21'b000011011011011001111};
                32'd1640 :tmp = {11'b0,21'b000011011011011100110};
                32'd1644 :tmp = {11'b0,21'b000011011011011101101};
                32'd1648 :tmp = {11'b0,21'b000011011011011111101};
                32'd1652 :tmp = {11'b0,21'b000011011011010000111};
                32'd1656 :tmp = {11'b0,21'b000011011011011111111};
                32'd1660 :tmp = {11'b0,21'b000011011011011101111};
                32'd1664 :tmp = {11'b0,21'b000011011111010111111};
                32'd1668 :tmp = {11'b0,21'b000011011111010000110};
                32'd1672 :tmp = {11'b0,21'b000011011111011011011};
                32'd1676 :tmp = {11'b0,21'b000011011111011001111};
                32'd1680 :tmp = {11'b0,21'b000011011111011100110};
                32'd1684 :tmp = {11'b0,21'b000011011111011101101};
                32'd1688 :tmp = {11'b0,21'b000011011111011111101};
                32'd1692 :tmp = {11'b0,21'b000011011111010000111};
                32'd1696 :tmp = {11'b0,21'b000011011111011111111};
                32'd1700 :tmp = {11'b0,21'b000011011111011101111};
                32'd1704 :tmp = {11'b0,21'b000011000001110111111};
                32'd1708 :tmp = {11'b0,21'b000011000001110000110};
                32'd1712 :tmp = {11'b0,21'b000011000001111011011};
                32'd1716 :tmp = {11'b0,21'b000011000001111001111};
                32'd1720 :tmp = {11'b0,21'b000011000001111100110};
                32'd1724 :tmp = {11'b0,21'b000011000001111101101};
                32'd1728 :tmp = {11'b0,21'b000011000001111111101};
                32'd1732 :tmp = {11'b0,21'b000011000001110000111};
                32'd1736 :tmp = {11'b0,21'b000011000001111111111};
                32'd1740 :tmp = {11'b0,21'b000011000001111101111};
                32'd1744 :tmp = {11'b0,21'b000011011111110111111};
                32'd1748 :tmp = {11'b0,21'b000011011111110000110};
                32'd1752 :tmp = {11'b0,21'b000011011111111011011};
                32'd1756 :tmp = {11'b0,21'b000011011111111001111};
                32'd1760 :tmp = {11'b0,21'b000011011111111100110};
                32'd1764 :tmp = {11'b0,21'b000011011111111101101};
                32'd1768 :tmp = {11'b0,21'b000011011111111111101};
                32'd1772 :tmp = {11'b0,21'b000011011111110000111};
                32'd1776 :tmp = {11'b0,21'b000011011111111111111};
                32'd1780 :tmp = {11'b0,21'b000011011111111101111};
                32'd1784 :tmp = {11'b0,21'b000011011011110111111};
                32'd1788 :tmp = {11'b0,21'b000011011011110000110};
                32'd1792 :tmp = {11'b0,21'b000011011011111011011};
                32'd1796 :tmp = {11'b0,21'b000011011011111001111};
                32'd1800 :tmp = {11'b0,21'b000011011011111100110};
                32'd1804 :tmp = {11'b0,21'b000011011011111101101};
                32'd1808 :tmp = {11'b0,21'b000011011011111111101};
                32'd1812 :tmp = {11'b0,21'b000011011011110000111};
                32'd1816 :tmp = {11'b0,21'b000011011011111111111};
                32'd1820 :tmp = {11'b0,21'b000011011011111101111};
                32'd1824 :tmp = {11'b0,21'b101101101111110111111};
                32'd1828 :tmp = {11'b0,21'b101101101111110000110};
                32'd1832 :tmp = {11'b0,21'b101101101111111011011};
                32'd1836 :tmp = {11'b0,21'b101101101111111001111};
                32'd1840 :tmp = {11'b0,21'b101101101111111100110};
                32'd1844 :tmp = {11'b0,21'b101101101111111101101};
                32'd1848 :tmp = {11'b0,21'b101101101111111111101};
                32'd1852 :tmp = {11'b0,21'b101101101111110000111};
                32'd1856 :tmp = {11'b0,21'b101101101111111111111};
                32'd1860 :tmp = {11'b0,21'b101101101111111101111};
                32'd1864 :tmp = {11'b0,21'b101101100001100111111};
                32'd1868 :tmp = {11'b0,21'b101101100001100000110};
                32'd1872 :tmp = {11'b0,21'b101101100001101011011};
                32'd1876 :tmp = {11'b0,21'b101101100001101001111};
                32'd1880 :tmp = {11'b0,21'b101101100001101100110};
                32'd1884 :tmp = {11'b0,21'b101101100001101101101};
                32'd1888 :tmp = {11'b0,21'b101101100001101111101};
                32'd1892 :tmp = {11'b0,21'b101101100001100000111};
                32'd1896 :tmp = {11'b0,21'b101101100001101111111};
                32'd1900 :tmp = {11'b0,21'b101101100001101101111};
                32'd1904 :tmp = {11'b0,21'b101101110110110111111};
                32'd1908 :tmp = {11'b0,21'b101101110110110000110};
                32'd1912 :tmp = {11'b0,21'b101101110110111011011};
                32'd1916 :tmp = {11'b0,21'b101101110110111001111};
                32'd1920 :tmp = {11'b0,21'b101101110110111100110};
                32'd1924 :tmp = {11'b0,21'b101101110110111101101};
                32'd1928 :tmp = {11'b0,21'b101101110110111111101};
                32'd1932 :tmp = {11'b0,21'b101101110110110000111};
                32'd1936 :tmp = {11'b0,21'b101101110110111111111};
                32'd1940 :tmp = {11'b0,21'b101101110110111101111};
                32'd1944 :tmp = {11'b0,21'b101101110011110111111};
                32'd1948 :tmp = {11'b0,21'b101101110011110000110};
                32'd1952 :tmp = {11'b0,21'b101101110011111011011};
                32'd1956 :tmp = {11'b0,21'b101101110011111001111};
                32'd1960 :tmp = {11'b0,21'b101101110011111100110};
                32'd1964 :tmp = {11'b0,21'b101101110011111101101};
                32'd1968 :tmp = {11'b0,21'b101101110011111111101};
                32'd1972 :tmp = {11'b0,21'b101101110011110000111};
                32'd1976 :tmp = {11'b0,21'b101101110011111111111};
                32'd1980 :tmp = {11'b0,21'b101101110011111101111};
                32'd1984 :tmp = {11'b0,21'b101101111001100111111};
                32'd1988 :tmp = {11'b0,21'b101101111001100000110};
                32'd1992 :tmp = {11'b0,21'b101101111001101011011};
                32'd1996 :tmp = {11'b0,21'b101101111001101001111};
                32'd2000 :tmp = {11'b0,21'b101101111001101100110};
                32'd2004 :tmp = {11'b0,21'b101101111001101101101};
                32'd2008 :tmp = {11'b0,21'b101101111001101111101};
                32'd2012 :tmp = {11'b0,21'b101101111001100000111};
                32'd2016 :tmp = {11'b0,21'b101101111001101111111};
                32'd2020 :tmp = {11'b0,21'b101101111001101101111};
                32'd2024 :tmp = {11'b0,21'b101101111011010111111};
                32'd2028 :tmp = {11'b0,21'b101101111011010000110};
                32'd2032 :tmp = {11'b0,21'b101101111011011011011};
                32'd2036 :tmp = {11'b0,21'b101101111011011001111};
                32'd2040 :tmp = {11'b0,21'b101101111011011100110};
                32'd2044 :tmp = {11'b0,21'b101101111011011101101};
                default : tmp = memory[address[9:2]];
            endcase end
            else tmp = 32'b0;

    always@ (posedge reset or posedge clk)
    if(reset)
        for (i = 0; i < 256; i = i + 1)
        memory[i] <= 32'h00000000;
    else begin 
        if(write_enable) begin
            if(Uart_send_trigger == 1'b1) Uart_send_trigger = 1'b0;
            case(address)
                32'h40000018 : begin UartWriteData <= writedata[7:0]; Uart_send_trigger <= 1'b1; end
                32'h40000014 : tubereg <= writedata[17:0];
                32'h4000000C : ledreg <= writedata[7:0];
                32'h40000000 : timer_TH <= writedata;
                32'h40000008 : timer_CON_W <= writedata[1:0];
                32'h40000020 : Uart_CON_W <= writedata[1:0];
                default : memory[address[9:2]] <= writedata;
            endcase 
            end
        end
    
    assign if_continue = timer_CON_R;
    Timer timer(clk,timer_CON_W,timer_TH,timer_CON_R,timer_TL);
    UART Uart(sysclk,Uart_state_trigger,Uart_Rx,UartWriteData,Uart_CON_W[1],Uart_CON_W[0],Uart_send_trigger,Uart_CON_R[0],Uart_CON_R[1],Uart_CON_R[2],Uart_Tx,UartReadData);
endmodule
